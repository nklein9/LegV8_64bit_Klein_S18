//Nicholas Klein
//Last Edit Feb 19, 2018
module programCounter();
	output PC;
	output PC4;
	input PS;
	input in;

endmodule
