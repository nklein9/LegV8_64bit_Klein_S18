module Mux64to1(a, s, out);
	//inputs and outputs
	input [63:0]a;
	input [5:0]s;
	output reg out;
	
	always @(*) begin
	case (s)
		6'b000000: out <= a[0];
		6'b000001: out <= a[1];
		6'b000010: out <= a[2];
		6'b000011: out <= a[3];
		6'b000100: out <= a[4];
		6'b000101: out <= a[5];
		6'b000110: out <= a[6];
		6'b000111: out <= a[7];
		6'b001000: out <= a[8];
		6'b001001: out <= a[9];
		6'b001010: out <= a[10];
		6'b001011: out <= a[11];
		6'b001100: out <= a[12];
		6'b001101: out <= a[13];
		6'b001110: out <= a[14];
		6'b001111: out <= a[15];
		6'b010000: out <= a[16];
		6'b010001: out <= a[17];
		6'b010010: out <= a[18];
		6'b010011: out <= a[19];
		6'b010100: out <= a[20];
		6'b010101: out <= a[21];
		6'b010110: out <= a[22];
		6'b010111: out <= a[23];
		6'b011000: out <= a[24];
		6'b011001: out <= a[25];
		6'b011010: out <= a[26];
		6'b011011: out <= a[27];
		6'b011100: out <= a[28];
		6'b011101: out <= a[29];
		6'b011110: out <= a[30];
		6'b011111: out <= a[31];
		6'b100000: out <= a[32];
		6'b100001: out <= a[33];
		6'b100010: out <= a[34];
		6'b100011: out <= a[35];
		6'b100100: out <= a[36];
		6'b100101: out <= a[37];
		6'b100110: out <= a[38];
		6'b100111: out <= a[39];
		6'b101000: out <= a[40];
		6'b101001: out <= a[41];
		6'b101010: out <= a[42];
		6'b101011: out <= a[43];
		6'b101100: out <= a[44];
		6'b101101: out <= a[45];
		6'b101110: out <= a[46];
		6'b101111: out <= a[47];
		6'b110000: out <= a[48];
		6'b110001: out <= a[49];
		6'b110010: out <= a[50];
		6'b110011: out <= a[51];
		6'b110100: out <= a[52];
		6'b110101: out <= a[53];
		6'b110110: out <= a[54];
		6'b110111: out <= a[55];
		6'b111000: out <= a[56];
		6'b111001: out <= a[57];
		6'b111010: out <= a[58];
		6'b111011: out <= a[59];
		6'b111100: out <= a[60];
		6'b111101: out <= a[61];
		6'b111110: out <= a[62];
		6'b111111: out <= a[63];
		
		default: out <= a[0];
	endcase
	end
endmodule
