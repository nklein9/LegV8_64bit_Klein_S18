//Nicholas Klein
//Last Edit Feb 19, 2018
module instructionRegister(out, in);
	output [31:0] out;
	input [31:0] in;

endmodule
